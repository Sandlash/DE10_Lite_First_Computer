// NiosII_esercitazione.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module NiosII_esercitazione (
		input  wire        clk_clk,            //         clk.clk
		output wire [7:0]  hex3_hex0_export,   //   hex3_hex0.export
		output wire [31:0] hex5_hex4_export,   //   hex5_hex4.export
		output wire [9:0]  leds_export,        //        leds.export
		input  wire [1:0]  push_button_export, // push_button.export
		input  wire        reset_reset_n,      //       reset.reset_n
		input  wire [9:0]  sliders_export      //     sliders.export
	);

	wire  [31:0] proc_data_master_readdata;                                   // mm_interconnect_0:proc_data_master_readdata -> proc:d_readdata
	wire         proc_data_master_waitrequest;                                // mm_interconnect_0:proc_data_master_waitrequest -> proc:d_waitrequest
	wire         proc_data_master_debugaccess;                                // proc:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:proc_data_master_debugaccess
	wire  [18:0] proc_data_master_address;                                    // proc:d_address -> mm_interconnect_0:proc_data_master_address
	wire   [3:0] proc_data_master_byteenable;                                 // proc:d_byteenable -> mm_interconnect_0:proc_data_master_byteenable
	wire         proc_data_master_read;                                       // proc:d_read -> mm_interconnect_0:proc_data_master_read
	wire         proc_data_master_write;                                      // proc:d_write -> mm_interconnect_0:proc_data_master_write
	wire  [31:0] proc_data_master_writedata;                                  // proc:d_writedata -> mm_interconnect_0:proc_data_master_writedata
	wire  [31:0] proc_instruction_master_readdata;                            // mm_interconnect_0:proc_instruction_master_readdata -> proc:i_readdata
	wire         proc_instruction_master_waitrequest;                         // mm_interconnect_0:proc_instruction_master_waitrequest -> proc:i_waitrequest
	wire  [18:0] proc_instruction_master_address;                             // proc:i_address -> mm_interconnect_0:proc_instruction_master_address
	wire         proc_instruction_master_read;                                // proc:i_read -> mm_interconnect_0:proc_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_proc_debug_mem_slave_readdata;             // proc:debug_mem_slave_readdata -> mm_interconnect_0:proc_debug_mem_slave_readdata
	wire         mm_interconnect_0_proc_debug_mem_slave_waitrequest;          // proc:debug_mem_slave_waitrequest -> mm_interconnect_0:proc_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_proc_debug_mem_slave_debugaccess;          // mm_interconnect_0:proc_debug_mem_slave_debugaccess -> proc:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_proc_debug_mem_slave_address;              // mm_interconnect_0:proc_debug_mem_slave_address -> proc:debug_mem_slave_address
	wire         mm_interconnect_0_proc_debug_mem_slave_read;                 // mm_interconnect_0:proc_debug_mem_slave_read -> proc:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_proc_debug_mem_slave_byteenable;           // mm_interconnect_0:proc_debug_mem_slave_byteenable -> proc:debug_mem_slave_byteenable
	wire         mm_interconnect_0_proc_debug_mem_slave_write;                // mm_interconnect_0:proc_debug_mem_slave_write -> proc:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_proc_debug_mem_slave_writedata;            // mm_interconnect_0:proc_debug_mem_slave_writedata -> proc:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_leds_s1_chipselect;                        // mm_interconnect_0:LEDs_s1_chipselect -> LEDs:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                          // LEDs:readdata -> mm_interconnect_0:LEDs_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                           // mm_interconnect_0:LEDs_s1_address -> LEDs:address
	wire         mm_interconnect_0_leds_s1_write;                             // mm_interconnect_0:LEDs_s1_write -> LEDs:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                         // mm_interconnect_0:LEDs_s1_writedata -> LEDs:writedata
	wire  [31:0] mm_interconnect_0_sliders_s1_readdata;                       // sliders:readdata -> mm_interconnect_0:sliders_s1_readdata
	wire   [1:0] mm_interconnect_0_sliders_s1_address;                        // mm_interconnect_0:sliders_s1_address -> sliders:address
	wire         mm_interconnect_0_hex3_hex0_s1_chipselect;                   // mm_interconnect_0:HEX3_HEX0_s1_chipselect -> HEX3_HEX0:chipselect
	wire  [31:0] mm_interconnect_0_hex3_hex0_s1_readdata;                     // HEX3_HEX0:readdata -> mm_interconnect_0:HEX3_HEX0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex3_hex0_s1_address;                      // mm_interconnect_0:HEX3_HEX0_s1_address -> HEX3_HEX0:address
	wire         mm_interconnect_0_hex3_hex0_s1_write;                        // mm_interconnect_0:HEX3_HEX0_s1_write -> HEX3_HEX0:write_n
	wire  [31:0] mm_interconnect_0_hex3_hex0_s1_writedata;                    // mm_interconnect_0:HEX3_HEX0_s1_writedata -> HEX3_HEX0:writedata
	wire         mm_interconnect_0_hex5_hex4_s1_chipselect;                   // mm_interconnect_0:HEX5_HEX4_s1_chipselect -> HEX5_HEX4:chipselect
	wire  [31:0] mm_interconnect_0_hex5_hex4_s1_readdata;                     // HEX5_HEX4:readdata -> mm_interconnect_0:HEX5_HEX4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex5_hex4_s1_address;                      // mm_interconnect_0:HEX5_HEX4_s1_address -> HEX5_HEX4:address
	wire         mm_interconnect_0_hex5_hex4_s1_write;                        // mm_interconnect_0:HEX5_HEX4_s1_write -> HEX5_HEX4:write_n
	wire  [31:0] mm_interconnect_0_hex5_hex4_s1_writedata;                    // mm_interconnect_0:HEX5_HEX4_s1_writedata -> HEX5_HEX4:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_watchdog_s1_chipselect;                    // mm_interconnect_0:watchdog_s1_chipselect -> watchdog:chipselect
	wire  [15:0] mm_interconnect_0_watchdog_s1_readdata;                      // watchdog:readdata -> mm_interconnect_0:watchdog_s1_readdata
	wire   [2:0] mm_interconnect_0_watchdog_s1_address;                       // mm_interconnect_0:watchdog_s1_address -> watchdog:address
	wire         mm_interconnect_0_watchdog_s1_write;                         // mm_interconnect_0:watchdog_s1_write -> watchdog:write_n
	wire  [15:0] mm_interconnect_0_watchdog_s1_writedata;                     // mm_interconnect_0:watchdog_s1_writedata -> watchdog:writedata
	wire         mm_interconnect_0_push_button_s1_chipselect;                 // mm_interconnect_0:push_button_s1_chipselect -> push_button:chipselect
	wire  [31:0] mm_interconnect_0_push_button_s1_readdata;                   // push_button:readdata -> mm_interconnect_0:push_button_s1_readdata
	wire   [1:0] mm_interconnect_0_push_button_s1_address;                    // mm_interconnect_0:push_button_s1_address -> push_button:address
	wire         mm_interconnect_0_push_button_s1_write;                      // mm_interconnect_0:push_button_s1_write -> push_button:write_n
	wire  [31:0] mm_interconnect_0_push_button_s1_writedata;                  // mm_interconnect_0:push_button_s1_writedata -> push_button:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s2_chipselect;            // mm_interconnect_0:onchip_memory2_0_s2_chipselect -> onchip_memory2_0:chipselect2
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s2_readdata;              // onchip_memory2_0:readdata2 -> mm_interconnect_0:onchip_memory2_0_s2_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_0_s2_address;               // mm_interconnect_0:onchip_memory2_0_s2_address -> onchip_memory2_0:address2
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s2_byteenable;            // mm_interconnect_0:onchip_memory2_0_s2_byteenable -> onchip_memory2_0:byteenable2
	wire         mm_interconnect_0_onchip_memory2_0_s2_write;                 // mm_interconnect_0:onchip_memory2_0_s2_write -> onchip_memory2_0:write2
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s2_writedata;             // mm_interconnect_0:onchip_memory2_0_s2_writedata -> onchip_memory2_0:writedata2
	wire         mm_interconnect_0_onchip_memory2_0_s2_clken;                 // mm_interconnect_0:onchip_memory2_0_s2_clken -> onchip_memory2_0:clken2
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // timer_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // push_button:irq -> irq_mapper:receiver2_irq
	wire  [31:0] proc_irq_irq;                                                // irq_mapper:sender_irq -> proc:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [HEX3_HEX0:reset_n, HEX5_HEX4:reset_n, LEDs:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:proc_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, proc:reset_n, push_button:reset_n, rst_translator:in_reset, sliders:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n, watchdog:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [onchip_memory2_0:reset_req, proc:reset_req, rst_translator:reset_req_in]
	wire         proc_debug_reset_request_reset;                              // proc:debug_reset_request -> rst_controller:reset_in1
	wire         watchdog_resetrequest_reset;                                 // watchdog:resetrequest -> rst_controller:reset_in2

	NiosII_esercitazione_HEX3_HEX0 hex3_hex0 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_hex3_hex0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex3_hex0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex3_hex0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex3_hex0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex3_hex0_s1_readdata),   //                    .readdata
		.out_port   (hex3_hex0_export)                           // external_connection.export
	);

	NiosII_esercitazione_HEX5_HEX4 hex5_hex4 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_hex5_hex4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex5_hex4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex5_hex4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex5_hex4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex5_hex4_s1_readdata),   //                    .readdata
		.out_port   (hex5_hex4_export)                           // external_connection.export
	);

	NiosII_esercitazione_LEDs leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	NiosII_esercitazione_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	NiosII_esercitazione_onchip_memory2_0 onchip_memory2_0 (
		.address     (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_0_onchip_memory2_0_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_onchip_memory2_0_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_onchip_memory2_0_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_onchip_memory2_0_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_onchip_memory2_0_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_onchip_memory2_0_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_onchip_memory2_0_s2_byteenable), //       .byteenable
		.clk         (clk_clk),                                          //   clk1.clk
		.reset       (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze      (1'b0)                                              // (terminated)
	);

	NiosII_esercitazione_proc proc (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (proc_data_master_address),                           //               data_master.address
		.d_byteenable                        (proc_data_master_byteenable),                        //                          .byteenable
		.d_read                              (proc_data_master_read),                              //                          .read
		.d_readdata                          (proc_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (proc_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (proc_data_master_write),                             //                          .write
		.d_writedata                         (proc_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (proc_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (proc_instruction_master_address),                    //        instruction_master.address
		.i_read                              (proc_instruction_master_read),                       //                          .read
		.i_readdata                          (proc_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (proc_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (proc_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (proc_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_proc_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_proc_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_proc_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_proc_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_proc_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_proc_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_proc_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_proc_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	NiosII_esercitazione_push_button push_button (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_push_button_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_push_button_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_push_button_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_push_button_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_push_button_s1_readdata),   //                    .readdata
		.in_port    (push_button_export),                          // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                     //                 irq.irq
	);

	NiosII_esercitazione_sliders sliders (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_sliders_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sliders_s1_readdata), //                    .readdata
		.in_port  (sliders_export)                         // external_connection.export
	);

	NiosII_esercitazione_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	NiosII_esercitazione_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	NiosII_esercitazione_watchdog watchdog (
		.clk          (clk_clk),                                  //          clk.clk
		.reset_n      (~rst_controller_reset_out_reset),          //        reset.reset_n
		.address      (mm_interconnect_0_watchdog_s1_address),    //           s1.address
		.writedata    (mm_interconnect_0_watchdog_s1_writedata),  //             .writedata
		.readdata     (mm_interconnect_0_watchdog_s1_readdata),   //             .readdata
		.chipselect   (mm_interconnect_0_watchdog_s1_chipselect), //             .chipselect
		.write_n      (~mm_interconnect_0_watchdog_s1_write),     //             .write_n
		.irq          (),                                         //          irq.irq
		.resetrequest (watchdog_resetrequest_reset)               // resetrequest.reset
	);

	NiosII_esercitazione_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                             (clk_clk),                                                     //                        clk_0_clk.clk
		.proc_reset_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                              // proc_reset_reset_bridge_in_reset.reset
		.proc_data_master_address                  (proc_data_master_address),                                    //                 proc_data_master.address
		.proc_data_master_waitrequest              (proc_data_master_waitrequest),                                //                                 .waitrequest
		.proc_data_master_byteenable               (proc_data_master_byteenable),                                 //                                 .byteenable
		.proc_data_master_read                     (proc_data_master_read),                                       //                                 .read
		.proc_data_master_readdata                 (proc_data_master_readdata),                                   //                                 .readdata
		.proc_data_master_write                    (proc_data_master_write),                                      //                                 .write
		.proc_data_master_writedata                (proc_data_master_writedata),                                  //                                 .writedata
		.proc_data_master_debugaccess              (proc_data_master_debugaccess),                                //                                 .debugaccess
		.proc_instruction_master_address           (proc_instruction_master_address),                             //          proc_instruction_master.address
		.proc_instruction_master_waitrequest       (proc_instruction_master_waitrequest),                         //                                 .waitrequest
		.proc_instruction_master_read              (proc_instruction_master_read),                                //                                 .read
		.proc_instruction_master_readdata          (proc_instruction_master_readdata),                            //                                 .readdata
		.HEX3_HEX0_s1_address                      (mm_interconnect_0_hex3_hex0_s1_address),                      //                     HEX3_HEX0_s1.address
		.HEX3_HEX0_s1_write                        (mm_interconnect_0_hex3_hex0_s1_write),                        //                                 .write
		.HEX3_HEX0_s1_readdata                     (mm_interconnect_0_hex3_hex0_s1_readdata),                     //                                 .readdata
		.HEX3_HEX0_s1_writedata                    (mm_interconnect_0_hex3_hex0_s1_writedata),                    //                                 .writedata
		.HEX3_HEX0_s1_chipselect                   (mm_interconnect_0_hex3_hex0_s1_chipselect),                   //                                 .chipselect
		.HEX5_HEX4_s1_address                      (mm_interconnect_0_hex5_hex4_s1_address),                      //                     HEX5_HEX4_s1.address
		.HEX5_HEX4_s1_write                        (mm_interconnect_0_hex5_hex4_s1_write),                        //                                 .write
		.HEX5_HEX4_s1_readdata                     (mm_interconnect_0_hex5_hex4_s1_readdata),                     //                                 .readdata
		.HEX5_HEX4_s1_writedata                    (mm_interconnect_0_hex5_hex4_s1_writedata),                    //                                 .writedata
		.HEX5_HEX4_s1_chipselect                   (mm_interconnect_0_hex5_hex4_s1_chipselect),                   //                                 .chipselect
		.jtag_uart_0_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //    jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                 .write
		.jtag_uart_0_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                 .read
		.jtag_uart_0_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                 .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                 .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                 .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                 .chipselect
		.LEDs_s1_address                           (mm_interconnect_0_leds_s1_address),                           //                          LEDs_s1.address
		.LEDs_s1_write                             (mm_interconnect_0_leds_s1_write),                             //                                 .write
		.LEDs_s1_readdata                          (mm_interconnect_0_leds_s1_readdata),                          //                                 .readdata
		.LEDs_s1_writedata                         (mm_interconnect_0_leds_s1_writedata),                         //                                 .writedata
		.LEDs_s1_chipselect                        (mm_interconnect_0_leds_s1_chipselect),                        //                                 .chipselect
		.onchip_memory2_0_s1_address               (mm_interconnect_0_onchip_memory2_0_s1_address),               //              onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                 (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                 .write
		.onchip_memory2_0_s1_readdata              (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                 .readdata
		.onchip_memory2_0_s1_writedata             (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                 .writedata
		.onchip_memory2_0_s1_byteenable            (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                 .byteenable
		.onchip_memory2_0_s1_chipselect            (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                 .chipselect
		.onchip_memory2_0_s1_clken                 (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                 .clken
		.onchip_memory2_0_s2_address               (mm_interconnect_0_onchip_memory2_0_s2_address),               //              onchip_memory2_0_s2.address
		.onchip_memory2_0_s2_write                 (mm_interconnect_0_onchip_memory2_0_s2_write),                 //                                 .write
		.onchip_memory2_0_s2_readdata              (mm_interconnect_0_onchip_memory2_0_s2_readdata),              //                                 .readdata
		.onchip_memory2_0_s2_writedata             (mm_interconnect_0_onchip_memory2_0_s2_writedata),             //                                 .writedata
		.onchip_memory2_0_s2_byteenable            (mm_interconnect_0_onchip_memory2_0_s2_byteenable),            //                                 .byteenable
		.onchip_memory2_0_s2_chipselect            (mm_interconnect_0_onchip_memory2_0_s2_chipselect),            //                                 .chipselect
		.onchip_memory2_0_s2_clken                 (mm_interconnect_0_onchip_memory2_0_s2_clken),                 //                                 .clken
		.proc_debug_mem_slave_address              (mm_interconnect_0_proc_debug_mem_slave_address),              //             proc_debug_mem_slave.address
		.proc_debug_mem_slave_write                (mm_interconnect_0_proc_debug_mem_slave_write),                //                                 .write
		.proc_debug_mem_slave_read                 (mm_interconnect_0_proc_debug_mem_slave_read),                 //                                 .read
		.proc_debug_mem_slave_readdata             (mm_interconnect_0_proc_debug_mem_slave_readdata),             //                                 .readdata
		.proc_debug_mem_slave_writedata            (mm_interconnect_0_proc_debug_mem_slave_writedata),            //                                 .writedata
		.proc_debug_mem_slave_byteenable           (mm_interconnect_0_proc_debug_mem_slave_byteenable),           //                                 .byteenable
		.proc_debug_mem_slave_waitrequest          (mm_interconnect_0_proc_debug_mem_slave_waitrequest),          //                                 .waitrequest
		.proc_debug_mem_slave_debugaccess          (mm_interconnect_0_proc_debug_mem_slave_debugaccess),          //                                 .debugaccess
		.push_button_s1_address                    (mm_interconnect_0_push_button_s1_address),                    //                   push_button_s1.address
		.push_button_s1_write                      (mm_interconnect_0_push_button_s1_write),                      //                                 .write
		.push_button_s1_readdata                   (mm_interconnect_0_push_button_s1_readdata),                   //                                 .readdata
		.push_button_s1_writedata                  (mm_interconnect_0_push_button_s1_writedata),                  //                                 .writedata
		.push_button_s1_chipselect                 (mm_interconnect_0_push_button_s1_chipselect),                 //                                 .chipselect
		.sliders_s1_address                        (mm_interconnect_0_sliders_s1_address),                        //                       sliders_s1.address
		.sliders_s1_readdata                       (mm_interconnect_0_sliders_s1_readdata),                       //                                 .readdata
		.sysid_qsys_0_control_slave_address        (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //       sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata       (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),       //                                 .readdata
		.timer_0_s1_address                        (mm_interconnect_0_timer_0_s1_address),                        //                       timer_0_s1.address
		.timer_0_s1_write                          (mm_interconnect_0_timer_0_s1_write),                          //                                 .write
		.timer_0_s1_readdata                       (mm_interconnect_0_timer_0_s1_readdata),                       //                                 .readdata
		.timer_0_s1_writedata                      (mm_interconnect_0_timer_0_s1_writedata),                      //                                 .writedata
		.timer_0_s1_chipselect                     (mm_interconnect_0_timer_0_s1_chipselect),                     //                                 .chipselect
		.watchdog_s1_address                       (mm_interconnect_0_watchdog_s1_address),                       //                      watchdog_s1.address
		.watchdog_s1_write                         (mm_interconnect_0_watchdog_s1_write),                         //                                 .write
		.watchdog_s1_readdata                      (mm_interconnect_0_watchdog_s1_readdata),                      //                                 .readdata
		.watchdog_s1_writedata                     (mm_interconnect_0_watchdog_s1_writedata),                     //                                 .writedata
		.watchdog_s1_chipselect                    (mm_interconnect_0_watchdog_s1_chipselect)                     //                                 .chipselect
	);

	NiosII_esercitazione_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (proc_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (proc_debug_reset_request_reset),     // reset_in1.reset
		.reset_in2      (watchdog_resetrequest_reset),        // reset_in2.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
